module not8bit(input [7:0] a,output [7:0] notout);

assign notout=~a;

endmodule